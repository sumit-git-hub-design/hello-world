module hello_world_tb;
 initial begin
   $display("Hello World");
   $finish;
 end
endmodule
